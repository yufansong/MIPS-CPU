`timescale 1ps/1ps

module InstructionMemory(Address, Instruction);
input [28:0] Address;
output [31:0] Instruction;

localparam ROM_SIZE = 1024;
reg [31:0] ROM[ROM_SIZE-1:0];
 
assign Instruction=(Address < ROM_SIZE)?ROM[Address]:32'b0;

integer i;
initial begin
for (i=0;i<ROM_SIZE;i=i+1) begin
            ROM[i] <= 32'h20100014;

// right
ROM[0] <= 32'h20100014;
ROM[1] <= 32'h20100014;
ROM[2] <= 32'h20100014;
ROM[3] <= 32'h20100014;
ROM[4] <= 32'h20050000;
ROM[5] <= 32'h3c051001;
ROM[5] <= 32'h20040001;
ROM[6] <= 32'h20090000;
ROM[7] <= 32'h200b0001;
ROM[8] <= 32'h200d0000;
ROM[9] <= 32'h200e0000;
ROM[10] <= 32'h01245020;
ROM[11] <= 32'h21490000;
ROM[12] <= 32'h01646020;
ROM[13] <= 32'h01846020;
ROM[14] <= 32'h01846020;
ROM[15] <= 32'h218b0000;
ROM[16] <= 32'h214d0000;
ROM[17] <= 32'h218e0000;
ROM[18] <= 32'h20840001;
ROM[19] <= 32'h1490fff6;
ROM[20] <= 32'h20100028;
ROM[21] <= 32'h01245020;
ROM[22] <= 32'h21490000;
ROM[23] <= 32'h01646020;
ROM[24] <= 32'h01846020;
ROM[25] <= 32'h01846020;
ROM[26] <= 32'h218b0000;
ROM[27] <= 32'h014c6820;
ROM[28] <= 32'h714d7002;
ROM[29] <= 32'h20840001;
ROM[30] <= 32'h1490fff6;
ROM[31] <= 32'h2010003c;
ROM[32] <= 32'h01245020;
ROM[33] <= 32'h21490000;
ROM[34] <= 32'h01646020;
ROM[35] <= 32'h01846020;
ROM[36] <= 32'h01846020;
ROM[37] <= 32'h218b0000;
ROM[38] <= 32'h714c6802;
ROM[39] <= 32'h718d7002;
// ROM[40] <= 32'h718d7002;
// ROM[41] <= 32'h718d7002;
// ROM[42] <= 32'h718d7002;
ROM[40] <= 32'h20840001;
ROM[41] <= 32'h1490fff6;

end
end
endmodule

// mul
// ROM[0] <= 32'h2004000a;
// ROM[1] <= 32'h2004000a;
// ROM[2] <= 32'h2004000a;
// ROM[3] <= 32'h2004000a;
// ROM[4] <= 32'h2005000d;
// ROM[5] <= 32'h70a43002;

//add a
// ROM[0] <= 32'h20090000;
// ROM[1] <= 32'h20090000;
// ROM[2] <= 32'h20090000;
// ROM[3] <= 32'h20090000;
// ROM[4] <= 32'h2010003c;
// ROM[5] <= 32'h20050000;
// ROM[6] <= 32'h3c050000;//ROM[6] <= 32'h3c051001;
// ROM[7] <= 32'h20040001;
// ROM[8] <= 32'haca90000;
// ROM[9] <= 32'h01245020;
// ROM[10] <= 32'h20a50004;
// ROM[11] <= 32'hacaa0000;
// ROM[12] <= 32'h20840001;
// ROM[13] <= 32'h21490000;
// ROM[14] <= 32'h1490fffa;


//original
// ROM[0] <= 32'b00001000000000000000000000000011;
// ROM[1] <= 32'b00001000000000000000000000101000;
// ROM[2] <= 32'b00001000000000000000000010010110;
// ROM[3] <= 32'b00001100000000000000000010010111;
// ROM[4] <= 32'b00100000000111010000000001000000;
// ROM[5] <= 32'b00111100000100000100000000000000;
// ROM[6] <= 32'b00100000000011000000000000000000;
// ROM[7] <= 32'b00111100000010011111111111111111;
// ROM[8] <= 32'b00100000000010011000000000000000;
// ROM[9] <= 32'b10101110000010010000000000000000;
// ROM[10] <= 32'b10101110000010010000000000000100;
// ROM[11] <= 32'b10101110000000000000000000001000;
// ROM[12] <= 32'b10101110000000000000000000001100;
// ROM[13] <= 32'b00100000000010010000000000000000;
// ROM[14] <= 32'b10101110000010010000000000010100;
// ROM[15] <= 32'b00100000000010010000000000000011;
// ROM[16] <= 32'b10101110000010010000000000100000;
// ROM[17] <= 32'b10001110000010100000000000100000;
// ROM[18] <= 32'b00110001010010010000000000001000;
// ROM[19] <= 32'b00010001001000001111111111111101;
// ROM[20] <= 32'b10001110000001010000000000011100;
// ROM[21] <= 32'b10001110000010100000000000100000;
// ROM[22] <= 32'b00110001010010010000000000001000;
// ROM[23] <= 32'b00010001001000001111111111111101;
// ROM[24] <= 32'b10001110000001100000000000011100;
// ROM[25] <= 32'b00100000000010010000000000000011;
// ROM[26] <= 32'b10101110000010010000000000001000;
// ROM[27] <= 32'b00100000101011010000000000000000;
// ROM[28] <= 32'b00100000110011100000000000000000;
// ROM[29] <= 32'b00010001101011100000000000000110;
// ROM[30] <= 32'b00000001101011100111100000101010;
// ROM[31] <= 32'b00010001111000000000000000000010;
// ROM[32] <= 32'b00000001110011010111000000100010;
// ROM[33] <= 32'b00001000000000000000000000011101;
// ROM[34] <= 32'b00000001101011100110100000100010;
// ROM[35] <= 32'b00001000000000000000000000011101;
// ROM[36] <= 32'b00100001110000110000000000000000;
// ROM[37] <= 32'b10101110000000110000000000001100;
// ROM[38] <= 32'b10101110000000110000000000011000;
// ROM[39] <= 32'b00001000000000000000000000010001;
// ROM[40] <= 32'b00100011101111011111111111111100;
// ROM[41] <= 32'b10101111101111110000000000000000;
// ROM[42] <= 32'b00111100000101111111111111111111;
// ROM[43] <= 32'b00100010111101111111111111111001;
// ROM[44] <= 32'b10001110000110000000000000001000;
// ROM[45] <= 32'b00000011000101111100000000100100;
// ROM[46] <= 32'b10101110000110000000000000001000;
// ROM[47] <= 32'b00010001100000000000000000000110;
// ROM[48] <= 32'b00100000000110010000000000000001;
// ROM[49] <= 32'b00010001100110010000000000001010;
// ROM[50] <= 32'b00100000000110010000000000000010;
// ROM[51] <= 32'b00010001100110010000000000001110;
// ROM[52] <= 32'b00100000000110010000000000000011;
// ROM[53] <= 32'b00010001100110010000000000010010;
// ROM[54] <= 32'b00000000000001011010011000000000;
// ROM[55] <= 32'b00000000000101001010011100000010;
// ROM[56] <= 32'b00001100000000000000000001001110;
// ROM[57] <= 32'b00100000111001110000100000000000;
// ROM[58] <= 32'b00100000000011000000000000000001;
// ROM[59] <= 32'b00001000000000000000000010001101;
// ROM[60] <= 32'b00000000000001011010011100000000;
// ROM[61] <= 32'b00000000000101001010011100000010;
// ROM[62] <= 32'b00001100000000000000000001001110;
// ROM[63] <= 32'b00100000111001110000010000000000;
// ROM[64] <= 32'b00100000000011000000000000000010;
// ROM[65] <= 32'b00001000000000000000000010001101;
// ROM[66] <= 32'b00000000000001101010011000000000;
// ROM[67] <= 32'b00000000000101001010011100000010;
// ROM[68] <= 32'b00001100000000000000000001001110;
// ROM[69] <= 32'b00100000111001110000001000000000;
// ROM[70] <= 32'b00100000000011000000000000000011;
// ROM[71] <= 32'b00001000000000000000000010001101;
// ROM[72] <= 32'b00000000000001101010011100000000;
// ROM[73] <= 32'b00000000000101001010011100000010;
// ROM[74] <= 32'b00001100000000000000000001001110;
// ROM[75] <= 32'b00100000111001110000000100000000;
// ROM[76] <= 32'b00100000000011000000000000000000;
// ROM[77] <= 32'b00001000000000000000000010001101;
// ROM[78] <= 32'b00100010100101111111111111110001;
// ROM[79] <= 32'b00010010111000000000000000011101;
// ROM[80] <= 32'b00100010100101111111111111110010;
// ROM[81] <= 32'b00010010111000000000000000011101;
// ROM[82] <= 32'b00100010100101111111111111110011;
// ROM[83] <= 32'b00010010111000000000000000011101;
// ROM[84] <= 32'b00100010100101111111111111110100;
// ROM[85] <= 32'b00010010111000000000000000011101;
// ROM[86] <= 32'b00100010100101111111111111110101;
// ROM[87] <= 32'b00010010111000000000000000011101;
// ROM[88] <= 32'b00100010100101111111111111110110;
// ROM[89] <= 32'b00010010111000000000000000011101;
// ROM[90] <= 32'b00100010100101111111111111110111;
// ROM[91] <= 32'b00010010111000000000000000011101;
// ROM[92] <= 32'b00100010100101111111111111111000;
// ROM[93] <= 32'b00010010111000000000000000011101;
// ROM[94] <= 32'b00100010100101111111111111111001;
// ROM[95] <= 32'b00010010111000000000000000011101;
// ROM[96] <= 32'b00100010100101111111111111111010;
// ROM[97] <= 32'b00010010111000000000000000011101;
// ROM[98] <= 32'b00100010100101111111111111111011;
// ROM[99] <= 32'b00010010111000000000000000011101;
// ROM[100] <= 32'b00100010100101111111111111111100;
// ROM[101] <= 32'b00010010111000000000000000011101;
// ROM[102] <= 32'b00100010100101111111111111111101;
// ROM[103] <= 32'b00010010111000000000000000011101;
// ROM[104] <= 32'b00100010100101111111111111111110;
// ROM[105] <= 32'b00010010111000000000000000011101;
// ROM[106] <= 32'b00100010100101111111111111111111;
// ROM[107] <= 32'b00010010111000000000000000011101;
// ROM[108] <= 32'b00010010100000000000000000011110;
// ROM[109] <= 32'b00100000000001110000000010001110;
// ROM[110] <= 32'b00000011111000000000000000001000;
// ROM[111] <= 32'b00100000000001110000000010011110;
// ROM[112] <= 32'b00000011111000000000000000001000;
// ROM[113] <= 32'b00100000000001110000000001111010;
// ROM[114] <= 32'b00000011111000000000000000001000;
// ROM[115] <= 32'b00100000000001110000000010011100;
// ROM[116] <= 32'b00000011111000000000000000001000;
// ROM[117] <= 32'b00100000000001110000000000111110;
// ROM[118] <= 32'b00000011111000000000000000001000;
// ROM[119] <= 32'b00100000000001110000000011101110;
// ROM[120] <= 32'b00000011111000000000000000001000;
// ROM[121] <= 32'b00100000000001110000000011110110;
// ROM[122] <= 32'b00000011111000000000000000001000;
// ROM[123] <= 32'b00100000000001110000000011111110;
// ROM[124] <= 32'b00000011111000000000000000001000;
// ROM[125] <= 32'b00100000000001110000000011100000;
// ROM[126] <= 32'b00000011111000000000000000001000;
// ROM[127] <= 32'b00100000000001110000000010111110;
// ROM[128] <= 32'b00000011111000000000000000001000;
// ROM[129] <= 32'b00100000000001110000000010110110;
// ROM[130] <= 32'b00000011111000000000000000001000;
// ROM[131] <= 32'b00100000000001110000000001100110;
// ROM[132] <= 32'b00000011111000000000000000001000;
// ROM[133] <= 32'b00100000000001110000000011110010;
// ROM[134] <= 32'b00000011111000000000000000001000;
// ROM[135] <= 32'b00100000000001110000000011011010;
// ROM[136] <= 32'b00000011111000000000000000001000;
// ROM[137] <= 32'b00100000000001110000000001100000;
// ROM[138] <= 32'b00000011111000000000000000001000;
// ROM[139] <= 32'b00100000000001110000000011111100;
// ROM[140] <= 32'b00000011111000000000000000001000;
// ROM[141] <= 32'b10001111101111110000000000000000;
// ROM[142] <= 32'b00100011101111010000000000000100;
// ROM[143] <= 32'b10101110000001110000000000010100;
// ROM[144] <= 32'b10001110000101010000000000001000;
// ROM[145] <= 32'b00100000000101100000000000000010;
// ROM[146] <= 32'b00000010101101101010100000100101;
// ROM[147] <= 32'b10101110000101010000000000001000;
// ROM[148] <= 32'b00100011010110101111111111111100;
// ROM[149] <= 32'b00000011010000000000000000001000;
// ROM[150] <= 32'b00000011010000000000000000001000;
// ROM[151] <= 32'b00000000000111111111100001000000;
// ROM[152] <= 32'b00000000000111111111100001000010;
// ROM[153] <= 32'b00000011111000000000000000001000;