module ALU(A, B, ALUFun, Sign, Z, Zero);
    input [31:0] A;
    input [31:0] B;
    input [5:0] ALUFun;
    input Sign; 
    
    output Zero;
    output [31:0] Z;
    
    wire [31:0] BOp;
    wire V, N, Zero;
    wire [31:0] AriOutput, BitOutput, ShiOutput, ComOutput;
    wire [31:0] SLL, SLL1, SLL2, SLL3, SLL4;
    wire [31:0] SRL, SRL1, SRL2, SRL3, SRL4;
    wire [31:0] SRA, SRA1, SRA2, SRA3, SRA4;
    //算术运算及指示位 add addu 00 sub subu 01  mul 10
    assign BOp = ALUFun[0] ? ~B+1 : B;
    assign AriOutput = ALUFun[1]? A * B:
                       (ALUFun[0] ?(A + ~B + 1) : A + B);
    
    assign Zero = (A == B) ? 0 : 1;
    // assign Zero = (A == B) ? 1 : 0;
    assign V = (Sign && (A[31] == BOp[31]) && (A[31] != AriOutput[31]))? 1:0;
    assign N = Sign ? (ALUFun[0] && AriOutput[31]) : (ALUFun[0] && A < B);
    
    //位运�?
    assign BitOutput = (ALUFun[3:0] == 4'b1000) ? A&B:
                       (ALUFun[3:0] == 4'b1110) ? A|B:
                       (ALUFun[3:0] == 4'b0110) ? A^B:
                       (ALUFun[3:0] == 4'b0001) ? ~(A|B):
                       (ALUFun[3:0] == 4'b1010) ? A: 32'b0; 
    
    //移位运算
    assign SLL = (A[4:0] == 5'b00000) ? B:
                 (A[4:0] == 5'b00001) ? {B[30:0], 1'b0}:
                 (A[4:0] == 5'b00010) ? {B[29:0], 2'b0}:
                 (A[4:0] == 5'b00011) ? {B[28:0], 3'b0}:
                 (A[4:0] == 5'b00100) ? {B[27:0], 4'b0}:
                 (A[4:0] == 5'b00101) ? {B[26:0], 5'b0}:
                 (A[4:0] == 5'b00110) ? {B[25:0], 6'b0}:
                 (A[4:0] == 5'b00111) ? {B[24:0], 7'b0}:
                 (A[4:0] == 5'b01000) ? {B[23:0], 8'b0}:
                 (A[4:0] == 5'b01001) ? {B[22:0], 9'b0}:
                 (A[4:0] == 5'b01010) ? {B[21:0], 10'b0}:
                 (A[4:0] == 5'b01011) ? {B[20:0], 11'b0}:
                 (A[4:0] == 5'b01100) ? {B[19:0], 12'b0}:
                 (A[4:0] == 5'b01101) ? {B[18:0], 13'b0}:
                 (A[4:0] == 5'b01110) ? {B[17:0], 14'b0}:
                 (A[4:0] == 5'b01111) ? {B[16:0], 15'b0}:
                 (A[4:0] == 5'b10000) ? {B[15:0], 16'b0}:
                 (A[4:0] == 5'b10001) ? {B[14:0], 17'b0}:
                 (A[4:0] == 5'b10010) ? {B[13:0], 18'b0}:
                 (A[4:0] == 5'b10011) ? {B[12:0], 19'b0}:
                 (A[4:0] == 5'b10100) ? {B[11:0], 20'b0}:
                 (A[4:0] == 5'b10101) ? {B[10:0], 21'b0}:
                 (A[4:0] == 5'b10110) ? {B[9:0], 22'b0}:
                 (A[4:0] == 5'b10111) ? {B[8:0], 23'b0}:
                 (A[4:0] == 5'b11000) ? {B[7:0], 24'b0}:
                 (A[4:0] == 5'b11001) ? {B[6:0], 25'b0}:
                 (A[4:0] == 5'b11010) ? {B[5:0], 26'b0}:
                 (A[4:0] == 5'b11011) ? {B[4:0], 27'b0}:
                 (A[4:0] == 5'b11100) ? {B[3:0], 28'b0}:
                 (A[4:0] == 5'b11101) ? {B[2:0], 29'b0}:
                 (A[4:0] == 5'b11110) ? {B[1:0], 30'b0}:
                 {B[0],31'b0};
    
    assign SRL = (A[4:0] == 5'b00000) ? B:
                 (A[4:0] == 5'b00001) ? {1'b0, B[31:1]}:
                 (A[4:0] == 5'b00010) ? {2'b0, B[31:2]}:
                 (A[4:0] == 5'b00011) ? {3'b0, B[31:3]}:
                 (A[4:0] == 5'b00100) ? {4'b0, B[31:4]}:
                 (A[4:0] == 5'b00101) ? {5'b0, B[31:5]}:
                 (A[4:0] == 5'b00110) ? {6'b0, B[31:6]}:
                 (A[4:0] == 5'b00111) ? {7'b0, B[31:7]}:
                 (A[4:0] == 5'b01000) ? {8'b0, B[31:8]}:
                 (A[4:0] == 5'b01001) ? {9'b0, B[31:9]}:
                 (A[4:0] == 5'b01010) ? {10'b0, B[31:10]}:
                 (A[4:0] == 5'b01011) ? {11'b0, B[31:11]}:
                 (A[4:0] == 5'b01100) ? {12'b0, B[31:12]}:
                 (A[4:0] == 5'b01101) ? {13'b0, B[31:13]}:
                 (A[4:0] == 5'b01110) ? {14'b0, B[31:14]}:
                 (A[4:0] == 5'b01111) ? {15'b0, B[31:15]}:
                 (A[4:0] == 5'b10000) ? {16'b0, B[31:16]}:
                 (A[4:0] == 5'b10001) ? {17'b0, B[31:17]}:
                 (A[4:0] == 5'b10010) ? {18'b0, B[31:18]}:
                 (A[4:0] == 5'b10011) ? {19'b0, B[31:19]}:
                 (A[4:0] == 5'b10100) ? {20'b0, B[31:20]}:
                 (A[4:0] == 5'b10101) ? {21'b0, B[31:21]}:
                 (A[4:0] == 5'b10110) ? {22'b0, B[31:22]}:
                 (A[4:0] == 5'b10111) ? {23'b0, B[31:23]}:
                 (A[4:0] == 5'b11000) ? {24'b0, B[31:24]}:
                 (A[4:0] == 5'b11001) ? {25'b0, B[31:25]}:
                 (A[4:0] == 5'b11010) ? {26'b0, B[31:26]}:
                 (A[4:0] == 5'b11011) ? {27'b0, B[31:27]}:
                 (A[4:0] == 5'b11100) ? {28'b0, B[31:28]}:
                 (A[4:0] == 5'b11101) ? {29'b0, B[31:29]}:
                 (A[4:0] == 5'b11110) ? {30'b0, B[31:30]}:
                 {31'b0, B[31]};
    
    assign SRA = (A[4:0] == 5'b00000) ? B:
                 (A[4:0] == 5'b00001) ? {B[31], B[31:1]}:
                 (A[4:0] == 5'b00010) ? {{2{B[31]}}, B[31:2]}:
                 (A[4:0] == 5'b00011) ? {{3{B[31]}}, B[31:3]}:
                 (A[4:0] == 5'b00100) ? {{4{B[31]}}, B[31:4]}:
                 (A[4:0] == 5'b00101) ? {{5{B[31]}}, B[31:5]}:
                 (A[4:0] == 5'b00110) ? {{6{B[31]}}, B[31:6]}:
                 (A[4:0] == 5'b00111) ? {{7{B[31]}}, B[31:7]}:
                 (A[4:0] == 5'b01000) ? {{8{B[31]}}, B[31:8]}:
                 (A[4:0] == 5'b01001) ? {{9{B[31]}}, B[31:9]}:
                 (A[4:0] == 5'b01010) ? {{10{B[31]}}, B[31:10]}:
                 (A[4:0] == 5'b01011) ? {{11{B[31]}}, B[31:11]}:
                 (A[4:0] == 5'b01100) ? {{12{B[31]}}, B[31:12]}:
                 (A[4:0] == 5'b01101) ? {{13{B[31]}}, B[31:13]}:
                 (A[4:0] == 5'b01110) ? {{14{B[31]}}, B[31:14]}:
                 (A[4:0] == 5'b01111) ? {{15{B[31]}}, B[31:15]}:
                 (A[4:0] == 5'b10000) ? {{16{B[31]}}, B[31:16]}:
                 (A[4:0] == 5'b10001) ? {{17{B[31]}}, B[31:17]}:
                 (A[4:0] == 5'b10010) ? {{18{B[31]}}, B[31:18]}:
                 (A[4:0] == 5'b10011) ? {{19{B[31]}}, B[31:19]}:
                 (A[4:0] == 5'b10100) ? {{20{B[31]}}, B[31:20]}:
                 (A[4:0] == 5'b10101) ? {{21{B[31]}}, B[31:21]}:
                 (A[4:0] == 5'b10110) ? {{22{B[31]}}, B[31:22]}:
                 (A[4:0] == 5'b10111) ? {{23{B[31]}}, B[31:23]}:
                 (A[4:0] == 5'b11000) ? {{24{B[31]}}, B[31:24]}:
                 (A[4:0] == 5'b11001) ? {{25{B[31]}}, B[31:25]}:
                 (A[4:0] == 5'b11010) ? {{26{B[31]}}, B[31:26]}:
                 (A[4:0] == 5'b11011) ? {{27{B[31]}}, B[31:27]}:
                 (A[4:0] == 5'b11100) ? {{28{B[31]}}, B[31:28]}:
                 (A[4:0] == 5'b11101) ? {{29{B[31]}}, B[31:29]}:
                 (A[4:0] == 5'b11110) ? {{30{B[31]}}, B[31:30]}:
                 {{31{B[31]}}, B[31]};
                 
    
    assign ShiOutput = (ALUFun[1:0] == 2'b00) ? SLL :
                       (ALUFun[1:0] == 2'b01) ? SRL :
                       (ALUFun[1:0] == 2'b11) ? SRA : 32'b0;
                       
    //关系运算
    assign ComOutput = (ALUFun[3:1] == 3'b001) ? {31'b0, Zero}:
                       (ALUFun[3:1] == 3'b000) ? {31'b0, ~Zero}:
                       (ALUFun[3:1] == 3'b010) ? {31'b0, N}:
                       (ALUFun[3:1] == 3'b110) ? {31'b0, (Sign&A[31])|(A==0)}:
                       (ALUFun[3:1] == 3'b101) ? {31'b0, Sign&A[31]}:
                       (ALUFun[3:1] == 3'b111) ? {31'b0, ~((Sign&A[31])|(A==0))}:32'b0;
   
   
    assign Z = (ALUFun[5:4] == 2'b00) ? AriOutput:
               (ALUFun[5:4] == 2'b01) ? BitOutput:
               (ALUFun[5:4] == 2'b10) ? ShiOutput:
               (ALUFun[5:4] == 2'b11) ? ComOutput: 32'b0;

endmodule